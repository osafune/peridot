-- pwm_control_core.vhd

-- Generated using ACDS version 13.1 162 at 2014.06.24.16:18:00

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pwm_control_core is
	port (
		clk_clk         : in  std_logic                    := '0'; --      clk.clk
		reset_reset_n   : in  std_logic                    := '0'; --    reset.reset_n
		pwm_data_export : out std_logic_vector(7 downto 0);        -- pwm_data.export
		scif_sclk       : in  std_logic                    := '0'; --     scif.sclk
		scif_txd        : in  std_logic                    := '0'; --         .txd
		scif_txr_n      : out std_logic;                           --         .txr_n
		scif_rxd        : out std_logic;                           --         .rxd
		scif_rxr_n      : in  std_logic                    := '0'  --         .rxr_n
	);
end entity pwm_control_core;

architecture rtl of pwm_control_core is
	component pwm_control_core_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component pwm_control_core_sysid;

	component pwm_control_core_pwmdata is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component pwm_control_core_pwmdata;

	component peridot_avalonmm_bridge is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			address       : out std_logic_vector(31 downto 0);                    -- address
			readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			read          : out std_logic;                                        -- read
			write         : out std_logic;                                        -- write
			byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			scif_sclk     : in  std_logic                     := 'X';             -- export
			scif_txd      : in  std_logic                     := 'X';             -- export
			scif_txr_n    : out std_logic;                                        -- export
			scif_rxd      : out std_logic;                                        -- export
			scif_rxr_n    : in  std_logic                     := 'X'              -- export
		);
	end component peridot_avalonmm_bridge;

	component pwm_control_core_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			peridot_bridge_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			peridot_bridge_avalon_master_address             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			peridot_bridge_avalon_master_waitrequest         : out std_logic;                                        -- waitrequest
			peridot_bridge_avalon_master_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			peridot_bridge_avalon_master_read                : in  std_logic                     := 'X';             -- read
			peridot_bridge_avalon_master_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			peridot_bridge_avalon_master_readdatavalid       : out std_logic;                                        -- readdatavalid
			peridot_bridge_avalon_master_write               : in  std_logic                     := 'X';             -- write
			peridot_bridge_avalon_master_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pwmdata_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pwmdata_s1_write                                 : out std_logic;                                        -- write
			pwmdata_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwmdata_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pwmdata_s1_chipselect                            : out std_logic;                                        -- chipselect
			sysid_control_slave_address                      : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component pwm_control_core_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal mm_interconnect_0_pwmdata_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwmdata_s1_writedata -> pwmdata:writedata
	signal mm_interconnect_0_pwmdata_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pwmdata_s1_address -> pwmdata:address
	signal mm_interconnect_0_pwmdata_s1_chipselect        : std_logic;                     -- mm_interconnect_0:pwmdata_s1_chipselect -> pwmdata:chipselect
	signal mm_interconnect_0_pwmdata_s1_write             : std_logic;                     -- mm_interconnect_0:pwmdata_s1_write -> mm_interconnect_0_pwmdata_s1_write:in
	signal mm_interconnect_0_pwmdata_s1_readdata          : std_logic_vector(31 downto 0); -- pwmdata:readdata -> mm_interconnect_0:pwmdata_s1_readdata
	signal peridot_bridge_avalon_master_waitrequest       : std_logic;                     -- mm_interconnect_0:peridot_bridge_avalon_master_waitrequest -> peridot_bridge:waitrequest
	signal peridot_bridge_avalon_master_writedata         : std_logic_vector(31 downto 0); -- peridot_bridge:writedata -> mm_interconnect_0:peridot_bridge_avalon_master_writedata
	signal peridot_bridge_avalon_master_address           : std_logic_vector(31 downto 0); -- peridot_bridge:address -> mm_interconnect_0:peridot_bridge_avalon_master_address
	signal peridot_bridge_avalon_master_write             : std_logic;                     -- peridot_bridge:write -> mm_interconnect_0:peridot_bridge_avalon_master_write
	signal peridot_bridge_avalon_master_read              : std_logic;                     -- peridot_bridge:read -> mm_interconnect_0:peridot_bridge_avalon_master_read
	signal peridot_bridge_avalon_master_readdata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:peridot_bridge_avalon_master_readdata -> peridot_bridge:readdata
	signal peridot_bridge_avalon_master_readdatavalid     : std_logic;                     -- mm_interconnect_0:peridot_bridge_avalon_master_readdatavalid -> peridot_bridge:readdatavalid
	signal peridot_bridge_avalon_master_byteenable        : std_logic_vector(3 downto 0);  -- peridot_bridge:byteenable -> mm_interconnect_0:peridot_bridge_avalon_master_byteenable
	signal mm_interconnect_0_sysid_control_slave_address  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_sysid_control_slave_readdata : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal rst_controller_reset_out_reset                 : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:peridot_bridge_reset_reset_bridge_in_reset_reset, peridot_bridge:reset, rst_controller_reset_out_reset:in]
	signal reset_reset_n_ports_inv                        : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_pwmdata_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_pwmdata_s1_write:inv -> pwmdata:write_n
	signal rst_controller_reset_out_reset_ports_inv       : std_logic;                     -- rst_controller_reset_out_reset:inv -> [pwmdata:reset_n, sysid:reset_n]

begin

	sysid : component pwm_control_core_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	pwmdata : component pwm_control_core_pwmdata
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_pwmdata_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwmdata_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwmdata_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwmdata_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwmdata_s1_readdata,        --                    .readdata
			out_port   => pwm_data_export                               -- external_connection.export
		);

	peridot_bridge : component peridot_avalonmm_bridge
		port map (
			clk           => clk_clk,                                    --         clock.clk
			reset         => rst_controller_reset_out_reset,             --         reset.reset
			address       => peridot_bridge_avalon_master_address,       -- avalon_master.address
			readdata      => peridot_bridge_avalon_master_readdata,      --              .readdata
			read          => peridot_bridge_avalon_master_read,          --              .read
			write         => peridot_bridge_avalon_master_write,         --              .write
			byteenable    => peridot_bridge_avalon_master_byteenable,    --              .byteenable
			writedata     => peridot_bridge_avalon_master_writedata,     --              .writedata
			waitrequest   => peridot_bridge_avalon_master_waitrequest,   --              .waitrequest
			readdatavalid => peridot_bridge_avalon_master_readdatavalid, --              .readdatavalid
			scif_sclk     => scif_sclk,                                  --   conduit_end.export
			scif_txd      => scif_txd,                                   --              .export
			scif_txr_n    => scif_txr_n,                                 --              .export
			scif_rxd      => scif_rxd,                                   --              .export
			scif_rxr_n    => scif_rxr_n                                  --              .export
		);

	mm_interconnect_0 : component pwm_control_core_mm_interconnect_0
		port map (
			clk_0_clk_clk                                    => clk_clk,                                        --                                  clk_0_clk.clk
			peridot_bridge_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                 -- peridot_bridge_reset_reset_bridge_in_reset.reset
			peridot_bridge_avalon_master_address             => peridot_bridge_avalon_master_address,           --               peridot_bridge_avalon_master.address
			peridot_bridge_avalon_master_waitrequest         => peridot_bridge_avalon_master_waitrequest,       --                                           .waitrequest
			peridot_bridge_avalon_master_byteenable          => peridot_bridge_avalon_master_byteenable,        --                                           .byteenable
			peridot_bridge_avalon_master_read                => peridot_bridge_avalon_master_read,              --                                           .read
			peridot_bridge_avalon_master_readdata            => peridot_bridge_avalon_master_readdata,          --                                           .readdata
			peridot_bridge_avalon_master_readdatavalid       => peridot_bridge_avalon_master_readdatavalid,     --                                           .readdatavalid
			peridot_bridge_avalon_master_write               => peridot_bridge_avalon_master_write,             --                                           .write
			peridot_bridge_avalon_master_writedata           => peridot_bridge_avalon_master_writedata,         --                                           .writedata
			pwmdata_s1_address                               => mm_interconnect_0_pwmdata_s1_address,           --                                 pwmdata_s1.address
			pwmdata_s1_write                                 => mm_interconnect_0_pwmdata_s1_write,             --                                           .write
			pwmdata_s1_readdata                              => mm_interconnect_0_pwmdata_s1_readdata,          --                                           .readdata
			pwmdata_s1_writedata                             => mm_interconnect_0_pwmdata_s1_writedata,         --                                           .writedata
			pwmdata_s1_chipselect                            => mm_interconnect_0_pwmdata_s1_chipselect,        --                                           .chipselect
			sysid_control_slave_address                      => mm_interconnect_0_sysid_control_slave_address,  --                        sysid_control_slave.address
			sysid_control_slave_readdata                     => mm_interconnect_0_sysid_control_slave_readdata  --                                           .readdata
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_pwmdata_s1_write_ports_inv <= not mm_interconnect_0_pwmdata_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of pwm_control_core
