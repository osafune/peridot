// cq_viola.v

// Generated using ACDS version 13.1 162 at 2014.06.24.16:32:28

`timescale 1 ps / 1 ps
module cq_viola (
		input  wire        core_clk,      //   core.clk
		input  wire        reset_reset_n, //  reset.reset_n
		input  wire        peri_clk,      //   peri.clk
		output wire        sysled_export, // sysled.export
		output wire [11:0] sdr_addr,      //    sdr.addr
		output wire [1:0]  sdr_ba,        //       .ba
		output wire        sdr_cas_n,     //       .cas_n
		output wire        sdr_cke,       //       .cke
		output wire        sdr_cs_n,      //       .cs_n
		inout  wire [15:0] sdr_dq,        //       .dq
		output wire [1:0]  sdr_dqm,       //       .dqm
		output wire        sdr_ras_n,     //       .ras_n
		output wire        sdr_we_n,      //       .we_n
		inout  wire [27:0] gpio_export,   //   gpio.export
		input  wire        epcs_MISO,     //   epcs.MISO
		output wire        epcs_MOSI,     //       .MOSI
		output wire        epcs_SCLK,     //       .SCLK
		output wire        epcs_SS_n,     //       .SS_n
		input  wire        scif_sclk,     //   scif.sclk
		input  wire        scif_txd,      //       .txd
		output wire        scif_txr_n,    //       .txr_n
		output wire        scif_rxd,      //       .rxd
		input  wire        scif_rxr_n     //       .rxr_n
	);

	wire         nios2_e_instruction_master_waitrequest;                    // mm_interconnect_0:nios2_e_instruction_master_waitrequest -> nios2_e:i_waitrequest
	wire  [27:0] nios2_e_instruction_master_address;                        // nios2_e:i_address -> mm_interconnect_0:nios2_e_instruction_master_address
	wire         nios2_e_instruction_master_read;                           // nios2_e:i_read -> mm_interconnect_0:nios2_e_instruction_master_read
	wire  [31:0] nios2_e_instruction_master_readdata;                       // mm_interconnect_0:nios2_e_instruction_master_readdata -> nios2_e:i_readdata
	wire         nios2_e_data_master_waitrequest;                           // mm_interconnect_0:nios2_e_data_master_waitrequest -> nios2_e:d_waitrequest
	wire  [31:0] nios2_e_data_master_writedata;                             // nios2_e:d_writedata -> mm_interconnect_0:nios2_e_data_master_writedata
	wire  [28:0] nios2_e_data_master_address;                               // nios2_e:d_address -> mm_interconnect_0:nios2_e_data_master_address
	wire         nios2_e_data_master_write;                                 // nios2_e:d_write -> mm_interconnect_0:nios2_e_data_master_write
	wire         nios2_e_data_master_read;                                  // nios2_e:d_read -> mm_interconnect_0:nios2_e_data_master_read
	wire  [31:0] nios2_e_data_master_readdata;                              // mm_interconnect_0:nios2_e_data_master_readdata -> nios2_e:d_readdata
	wire         nios2_e_data_master_debugaccess;                           // nios2_e:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_e_data_master_debugaccess
	wire   [3:0] nios2_e_data_master_byteenable;                            // nios2_e:d_byteenable -> mm_interconnect_0:nios2_e_data_master_byteenable
	wire         mm_interconnect_0_nios2_e_jtag_debug_module_waitrequest;   // nios2_e:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_e_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_e_jtag_debug_module_writedata;     // mm_interconnect_0:nios2_e_jtag_debug_module_writedata -> nios2_e:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_e_jtag_debug_module_address;       // mm_interconnect_0:nios2_e_jtag_debug_module_address -> nios2_e:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_e_jtag_debug_module_write;         // mm_interconnect_0:nios2_e_jtag_debug_module_write -> nios2_e:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_e_jtag_debug_module_read;          // mm_interconnect_0:nios2_e_jtag_debug_module_read -> nios2_e:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_e_jtag_debug_module_readdata;      // nios2_e:jtag_debug_module_readdata -> mm_interconnect_0:nios2_e_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_e_jtag_debug_module_debugaccess;   // mm_interconnect_0:nios2_e_jtag_debug_module_debugaccess -> nios2_e:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_e_jtag_debug_module_byteenable;    // mm_interconnect_0:nios2_e_jtag_debug_module_byteenable -> nios2_e:jtag_debug_module_byteenable
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire  [31:0] mm_interconnect_0_ipl_memory_s1_writedata;                 // mm_interconnect_0:ipl_memory_s1_writedata -> ipl_memory:writedata
	wire  [11:0] mm_interconnect_0_ipl_memory_s1_address;                   // mm_interconnect_0:ipl_memory_s1_address -> ipl_memory:address
	wire         mm_interconnect_0_ipl_memory_s1_chipselect;                // mm_interconnect_0:ipl_memory_s1_chipselect -> ipl_memory:chipselect
	wire         mm_interconnect_0_ipl_memory_s1_clken;                     // mm_interconnect_0:ipl_memory_s1_clken -> ipl_memory:clken
	wire         mm_interconnect_0_ipl_memory_s1_write;                     // mm_interconnect_0:ipl_memory_s1_write -> ipl_memory:write
	wire  [31:0] mm_interconnect_0_ipl_memory_s1_readdata;                  // ipl_memory:readdata -> mm_interconnect_0:ipl_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_ipl_memory_s1_byteenable;                // mm_interconnect_0:ipl_memory_s1_byteenable -> ipl_memory:byteenable
	wire         mm_interconnect_0_peripherals_bridge_s0_waitrequest;       // peripherals_bridge:s0_waitrequest -> mm_interconnect_0:peripherals_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_peripherals_bridge_s0_burstcount;        // mm_interconnect_0:peripherals_bridge_s0_burstcount -> peripherals_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_peripherals_bridge_s0_writedata;         // mm_interconnect_0:peripherals_bridge_s0_writedata -> peripherals_bridge:s0_writedata
	wire  [15:0] mm_interconnect_0_peripherals_bridge_s0_address;           // mm_interconnect_0:peripherals_bridge_s0_address -> peripherals_bridge:s0_address
	wire         mm_interconnect_0_peripherals_bridge_s0_write;             // mm_interconnect_0:peripherals_bridge_s0_write -> peripherals_bridge:s0_write
	wire         mm_interconnect_0_peripherals_bridge_s0_read;              // mm_interconnect_0:peripherals_bridge_s0_read -> peripherals_bridge:s0_read
	wire  [31:0] mm_interconnect_0_peripherals_bridge_s0_readdata;          // peripherals_bridge:s0_readdata -> mm_interconnect_0:peripherals_bridge_s0_readdata
	wire         mm_interconnect_0_peripherals_bridge_s0_debugaccess;       // mm_interconnect_0:peripherals_bridge_s0_debugaccess -> peripherals_bridge:s0_debugaccess
	wire         mm_interconnect_0_peripherals_bridge_s0_readdatavalid;     // peripherals_bridge:s0_readdatavalid -> mm_interconnect_0:peripherals_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_peripherals_bridge_s0_byteenable;        // mm_interconnect_0:peripherals_bridge_s0_byteenable -> peripherals_bridge:s0_byteenable
	wire         peridot_bridge_avalon_master_waitrequest;                  // mm_interconnect_0:peridot_bridge_avalon_master_waitrequest -> peridot_bridge:waitrequest
	wire  [31:0] peridot_bridge_avalon_master_writedata;                    // peridot_bridge:writedata -> mm_interconnect_0:peridot_bridge_avalon_master_writedata
	wire  [31:0] peridot_bridge_avalon_master_address;                      // peridot_bridge:address -> mm_interconnect_0:peridot_bridge_avalon_master_address
	wire         peridot_bridge_avalon_master_write;                        // peridot_bridge:write -> mm_interconnect_0:peridot_bridge_avalon_master_write
	wire         peridot_bridge_avalon_master_read;                         // peridot_bridge:read -> mm_interconnect_0:peridot_bridge_avalon_master_read
	wire  [31:0] peridot_bridge_avalon_master_readdata;                     // mm_interconnect_0:peridot_bridge_avalon_master_readdata -> peridot_bridge:readdata
	wire         peridot_bridge_avalon_master_readdatavalid;                // mm_interconnect_0:peridot_bridge_avalon_master_readdatavalid -> peridot_bridge:readdatavalid
	wire   [3:0] peridot_bridge_avalon_master_byteenable;                   // peridot_bridge:byteenable -> mm_interconnect_0:peridot_bridge_avalon_master_byteenable
	wire  [31:0] mm_interconnect_1_gpio_0_s1_writedata;                     // mm_interconnect_1:gpio_0_s1_writedata -> gpio_0:writedata
	wire   [1:0] mm_interconnect_1_gpio_0_s1_address;                       // mm_interconnect_1:gpio_0_s1_address -> gpio_0:address
	wire         mm_interconnect_1_gpio_0_s1_chipselect;                    // mm_interconnect_1:gpio_0_s1_chipselect -> gpio_0:chipselect
	wire         mm_interconnect_1_gpio_0_s1_write;                         // mm_interconnect_1:gpio_0_s1_write -> gpio_0:write_n
	wire  [31:0] mm_interconnect_1_gpio_0_s1_readdata;                      // gpio_0:readdata -> mm_interconnect_1:gpio_0_s1_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;             // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire  [15:0] mm_interconnect_1_epcs_spi_spi_control_port_writedata;     // mm_interconnect_1:epcs_spi_spi_control_port_writedata -> epcs_spi:data_from_cpu
	wire   [2:0] mm_interconnect_1_epcs_spi_spi_control_port_address;       // mm_interconnect_1:epcs_spi_spi_control_port_address -> epcs_spi:mem_addr
	wire         mm_interconnect_1_epcs_spi_spi_control_port_chipselect;    // mm_interconnect_1:epcs_spi_spi_control_port_chipselect -> epcs_spi:spi_select
	wire         mm_interconnect_1_epcs_spi_spi_control_port_write;         // mm_interconnect_1:epcs_spi_spi_control_port_write -> epcs_spi:write_n
	wire         mm_interconnect_1_epcs_spi_spi_control_port_read;          // mm_interconnect_1:epcs_spi_spi_control_port_read -> epcs_spi:read_n
	wire  [15:0] mm_interconnect_1_epcs_spi_spi_control_port_readdata;      // epcs_spi:data_to_cpu -> mm_interconnect_1:epcs_spi_spi_control_port_readdata
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                        // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire   [1:0] mm_interconnect_1_led_s1_address;                          // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_chipselect;                       // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire         mm_interconnect_1_led_s1_write;                            // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                         // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire  [15:0] mm_interconnect_1_systimer_s1_writedata;                   // mm_interconnect_1:systimer_s1_writedata -> systimer:writedata
	wire   [2:0] mm_interconnect_1_systimer_s1_address;                     // mm_interconnect_1:systimer_s1_address -> systimer:address
	wire         mm_interconnect_1_systimer_s1_chipselect;                  // mm_interconnect_1:systimer_s1_chipselect -> systimer:chipselect
	wire         mm_interconnect_1_systimer_s1_write;                       // mm_interconnect_1:systimer_s1_write -> systimer:write_n
	wire  [15:0] mm_interconnect_1_systimer_s1_readdata;                    // systimer:readdata -> mm_interconnect_1:systimer_s1_readdata
	wire   [0:0] peripherals_bridge_m0_burstcount;                          // peripherals_bridge:m0_burstcount -> mm_interconnect_1:peripherals_bridge_m0_burstcount
	wire         peripherals_bridge_m0_waitrequest;                         // mm_interconnect_1:peripherals_bridge_m0_waitrequest -> peripherals_bridge:m0_waitrequest
	wire  [15:0] peripherals_bridge_m0_address;                             // peripherals_bridge:m0_address -> mm_interconnect_1:peripherals_bridge_m0_address
	wire  [31:0] peripherals_bridge_m0_writedata;                           // peripherals_bridge:m0_writedata -> mm_interconnect_1:peripherals_bridge_m0_writedata
	wire         peripherals_bridge_m0_write;                               // peripherals_bridge:m0_write -> mm_interconnect_1:peripherals_bridge_m0_write
	wire         peripherals_bridge_m0_read;                                // peripherals_bridge:m0_read -> mm_interconnect_1:peripherals_bridge_m0_read
	wire  [31:0] peripherals_bridge_m0_readdata;                            // mm_interconnect_1:peripherals_bridge_m0_readdata -> peripherals_bridge:m0_readdata
	wire         peripherals_bridge_m0_debugaccess;                         // peripherals_bridge:m0_debugaccess -> mm_interconnect_1:peripherals_bridge_m0_debugaccess
	wire   [3:0] peripherals_bridge_m0_byteenable;                          // peripherals_bridge:m0_byteenable -> mm_interconnect_1:peripherals_bridge_m0_byteenable
	wire         peripherals_bridge_m0_readdatavalid;                       // mm_interconnect_1:peripherals_bridge_m0_readdatavalid -> peripherals_bridge:m0_readdatavalid
	wire  [31:0] nios2_e_d_irq_irq;                                         // irq_mapper:sender_irq -> nios2_e:d_irq
	wire         irq_mapper_receiver0_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                             // systimer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                  // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                         // jtag_uart:av_irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                  // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                         // epcs_spi:irq -> irq_synchronizer_002:receiver_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [ipl_memory:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, mm_interconnect_0:nios2_e_reset_n_reset_bridge_in_reset_reset, nios2_e:reset_n, peridot_bridge:reset, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [ipl_memory:reset_req, nios2_e:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [epcs_spi:reset_n, gpio_0:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:peripherals_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:peripherals_bridge_reset_reset_bridge_in_reset_reset, peripherals_bridge:reset, sysid:reset_n, systimer:reset_n]

	cq_viola_nios2_e nios2_e (
		.clk                                   (core_clk),                                                //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                         //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                             (nios2_e_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_e_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_e_data_master_read),                                //                          .read
		.d_readdata                            (nios2_e_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_e_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_e_data_master_write),                               //                          .write
		.d_writedata                           (nios2_e_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_e_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_e_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_e_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_e_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_e_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_e_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                        //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_e_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_e_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_e_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_e_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_e_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_e_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_e_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_e_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                         // custom_instruction_master.readra
	);

	cq_viola_jtag_uart jtag_uart (
		.clk            (peri_clk),                                                  //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_001_receiver_irq)                          //               irq.irq
	);

	cq_viola_ipl_memory ipl_memory (
		.clk        (core_clk),                                   //   clk1.clk
		.address    (mm_interconnect_0_ipl_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ipl_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ipl_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ipl_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ipl_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ipl_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ipl_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	cq_viola_sysid sysid (
		.clock    (peri_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	cq_viola_systimer systimer (
		.clk        (peri_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.address    (mm_interconnect_1_systimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_systimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_systimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_systimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_systimer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)             //   irq.irq
	);

	cq_viola_led led (
		.clk        (peri_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (sysled_export)                        // external_connection.export
	);

	cq_viola_sdram sdram (
		.clk            (core_clk),                                 //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdr_addr),                                 //  wire.export
		.zs_ba          (sdr_ba),                                   //      .export
		.zs_cas_n       (sdr_cas_n),                                //      .export
		.zs_cke         (sdr_cke),                                  //      .export
		.zs_cs_n        (sdr_cs_n),                                 //      .export
		.zs_dq          (sdr_dq),                                   //      .export
		.zs_dqm         (sdr_dqm),                                  //      .export
		.zs_ras_n       (sdr_ras_n),                                //      .export
		.zs_we_n        (sdr_we_n)                                  //      .export
	);

	cq_viola_gpio_0 gpio_0 (
		.clk        (peri_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_gpio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_gpio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_gpio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_gpio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_gpio_0_s1_readdata),   //                    .readdata
		.bidir_port (gpio_export)                             // external_connection.export
	);

	cq_viola_epcs_spi epcs_spi (
		.clk           (peri_clk),                                               //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                    //            reset.reset_n
		.data_from_cpu (mm_interconnect_1_epcs_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_1_epcs_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_1_epcs_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_1_epcs_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_1_epcs_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_1_epcs_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_synchronizer_002_receiver_irq),                      //              irq.irq
		.MISO          (epcs_MISO),                                              //         external.export
		.MOSI          (epcs_MOSI),                                              //                 .export
		.SCLK          (epcs_SCLK),                                              //                 .export
		.SS_n          (epcs_SS_n)                                               //                 .export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (16),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) peripherals_bridge (
		.clk              (peri_clk),                                              //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),                    // reset.reset
		.s0_waitrequest   (mm_interconnect_0_peripherals_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_peripherals_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_peripherals_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_peripherals_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_peripherals_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_peripherals_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_peripherals_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_peripherals_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_peripherals_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_peripherals_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (peripherals_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (peripherals_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (peripherals_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (peripherals_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (peripherals_bridge_m0_writedata),                       //      .writedata
		.m0_address       (peripherals_bridge_m0_address),                         //      .address
		.m0_write         (peripherals_bridge_m0_write),                           //      .write
		.m0_read          (peripherals_bridge_m0_read),                            //      .read
		.m0_byteenable    (peripherals_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (peripherals_bridge_m0_debugaccess)                      //      .debugaccess
	);

	peridot_avalonmm_bridge peridot_bridge (
		.clk           (core_clk),                                   //         clock.clk
		.reset         (rst_controller_reset_out_reset),             //         reset.reset
		.address       (peridot_bridge_avalon_master_address),       // avalon_master.address
		.readdata      (peridot_bridge_avalon_master_readdata),      //              .readdata
		.read          (peridot_bridge_avalon_master_read),          //              .read
		.write         (peridot_bridge_avalon_master_write),         //              .write
		.byteenable    (peridot_bridge_avalon_master_byteenable),    //              .byteenable
		.writedata     (peridot_bridge_avalon_master_writedata),     //              .writedata
		.waitrequest   (peridot_bridge_avalon_master_waitrequest),   //              .waitrequest
		.readdatavalid (peridot_bridge_avalon_master_readdatavalid), //              .readdatavalid
		.scif_sclk     (scif_sclk),                                  //   conduit_end.export
		.scif_txd      (scif_txd),                                   //              .export
		.scif_txr_n    (scif_txr_n),                                 //              .export
		.scif_rxd      (scif_rxd),                                   //              .export
		.scif_rxr_n    (scif_rxr_n)                                  //              .export
	);

	cq_viola_mm_interconnect_0 mm_interconnect_0 (
		.clk_core_clk_clk                                     (core_clk),                                                //                                   clk_core_clk.clk
		.clk_peri_clk_clk                                     (peri_clk),                                                //                                   clk_peri_clk.clk
		.nios2_e_reset_n_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                          //          nios2_e_reset_n_reset_bridge_in_reset.reset
		.peripherals_bridge_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                      // peripherals_bridge_reset_reset_bridge_in_reset.reset
		.nios2_e_data_master_address                          (nios2_e_data_master_address),                             //                            nios2_e_data_master.address
		.nios2_e_data_master_waitrequest                      (nios2_e_data_master_waitrequest),                         //                                               .waitrequest
		.nios2_e_data_master_byteenable                       (nios2_e_data_master_byteenable),                          //                                               .byteenable
		.nios2_e_data_master_read                             (nios2_e_data_master_read),                                //                                               .read
		.nios2_e_data_master_readdata                         (nios2_e_data_master_readdata),                            //                                               .readdata
		.nios2_e_data_master_write                            (nios2_e_data_master_write),                               //                                               .write
		.nios2_e_data_master_writedata                        (nios2_e_data_master_writedata),                           //                                               .writedata
		.nios2_e_data_master_debugaccess                      (nios2_e_data_master_debugaccess),                         //                                               .debugaccess
		.nios2_e_instruction_master_address                   (nios2_e_instruction_master_address),                      //                     nios2_e_instruction_master.address
		.nios2_e_instruction_master_waitrequest               (nios2_e_instruction_master_waitrequest),                  //                                               .waitrequest
		.nios2_e_instruction_master_read                      (nios2_e_instruction_master_read),                         //                                               .read
		.nios2_e_instruction_master_readdata                  (nios2_e_instruction_master_readdata),                     //                                               .readdata
		.peridot_bridge_avalon_master_address                 (peridot_bridge_avalon_master_address),                    //                   peridot_bridge_avalon_master.address
		.peridot_bridge_avalon_master_waitrequest             (peridot_bridge_avalon_master_waitrequest),                //                                               .waitrequest
		.peridot_bridge_avalon_master_byteenable              (peridot_bridge_avalon_master_byteenable),                 //                                               .byteenable
		.peridot_bridge_avalon_master_read                    (peridot_bridge_avalon_master_read),                       //                                               .read
		.peridot_bridge_avalon_master_readdata                (peridot_bridge_avalon_master_readdata),                   //                                               .readdata
		.peridot_bridge_avalon_master_readdatavalid           (peridot_bridge_avalon_master_readdatavalid),              //                                               .readdatavalid
		.peridot_bridge_avalon_master_write                   (peridot_bridge_avalon_master_write),                      //                                               .write
		.peridot_bridge_avalon_master_writedata               (peridot_bridge_avalon_master_writedata),                  //                                               .writedata
		.ipl_memory_s1_address                                (mm_interconnect_0_ipl_memory_s1_address),                 //                                  ipl_memory_s1.address
		.ipl_memory_s1_write                                  (mm_interconnect_0_ipl_memory_s1_write),                   //                                               .write
		.ipl_memory_s1_readdata                               (mm_interconnect_0_ipl_memory_s1_readdata),                //                                               .readdata
		.ipl_memory_s1_writedata                              (mm_interconnect_0_ipl_memory_s1_writedata),               //                                               .writedata
		.ipl_memory_s1_byteenable                             (mm_interconnect_0_ipl_memory_s1_byteenable),              //                                               .byteenable
		.ipl_memory_s1_chipselect                             (mm_interconnect_0_ipl_memory_s1_chipselect),              //                                               .chipselect
		.ipl_memory_s1_clken                                  (mm_interconnect_0_ipl_memory_s1_clken),                   //                                               .clken
		.nios2_e_jtag_debug_module_address                    (mm_interconnect_0_nios2_e_jtag_debug_module_address),     //                      nios2_e_jtag_debug_module.address
		.nios2_e_jtag_debug_module_write                      (mm_interconnect_0_nios2_e_jtag_debug_module_write),       //                                               .write
		.nios2_e_jtag_debug_module_read                       (mm_interconnect_0_nios2_e_jtag_debug_module_read),        //                                               .read
		.nios2_e_jtag_debug_module_readdata                   (mm_interconnect_0_nios2_e_jtag_debug_module_readdata),    //                                               .readdata
		.nios2_e_jtag_debug_module_writedata                  (mm_interconnect_0_nios2_e_jtag_debug_module_writedata),   //                                               .writedata
		.nios2_e_jtag_debug_module_byteenable                 (mm_interconnect_0_nios2_e_jtag_debug_module_byteenable),  //                                               .byteenable
		.nios2_e_jtag_debug_module_waitrequest                (mm_interconnect_0_nios2_e_jtag_debug_module_waitrequest), //                                               .waitrequest
		.nios2_e_jtag_debug_module_debugaccess                (mm_interconnect_0_nios2_e_jtag_debug_module_debugaccess), //                                               .debugaccess
		.peripherals_bridge_s0_address                        (mm_interconnect_0_peripherals_bridge_s0_address),         //                          peripherals_bridge_s0.address
		.peripherals_bridge_s0_write                          (mm_interconnect_0_peripherals_bridge_s0_write),           //                                               .write
		.peripherals_bridge_s0_read                           (mm_interconnect_0_peripherals_bridge_s0_read),            //                                               .read
		.peripherals_bridge_s0_readdata                       (mm_interconnect_0_peripherals_bridge_s0_readdata),        //                                               .readdata
		.peripherals_bridge_s0_writedata                      (mm_interconnect_0_peripherals_bridge_s0_writedata),       //                                               .writedata
		.peripherals_bridge_s0_burstcount                     (mm_interconnect_0_peripherals_bridge_s0_burstcount),      //                                               .burstcount
		.peripherals_bridge_s0_byteenable                     (mm_interconnect_0_peripherals_bridge_s0_byteenable),      //                                               .byteenable
		.peripherals_bridge_s0_readdatavalid                  (mm_interconnect_0_peripherals_bridge_s0_readdatavalid),   //                                               .readdatavalid
		.peripherals_bridge_s0_waitrequest                    (mm_interconnect_0_peripherals_bridge_s0_waitrequest),     //                                               .waitrequest
		.peripherals_bridge_s0_debugaccess                    (mm_interconnect_0_peripherals_bridge_s0_debugaccess),     //                                               .debugaccess
		.sdram_s1_address                                     (mm_interconnect_0_sdram_s1_address),                      //                                       sdram_s1.address
		.sdram_s1_write                                       (mm_interconnect_0_sdram_s1_write),                        //                                               .write
		.sdram_s1_read                                        (mm_interconnect_0_sdram_s1_read),                         //                                               .read
		.sdram_s1_readdata                                    (mm_interconnect_0_sdram_s1_readdata),                     //                                               .readdata
		.sdram_s1_writedata                                   (mm_interconnect_0_sdram_s1_writedata),                    //                                               .writedata
		.sdram_s1_byteenable                                  (mm_interconnect_0_sdram_s1_byteenable),                   //                                               .byteenable
		.sdram_s1_readdatavalid                               (mm_interconnect_0_sdram_s1_readdatavalid),                //                                               .readdatavalid
		.sdram_s1_waitrequest                                 (mm_interconnect_0_sdram_s1_waitrequest),                  //                                               .waitrequest
		.sdram_s1_chipselect                                  (mm_interconnect_0_sdram_s1_chipselect)                    //                                               .chipselect
	);

	cq_viola_mm_interconnect_1 mm_interconnect_1 (
		.clk_peri_clk_clk                                     (peri_clk),                                                  //                                   clk_peri_clk.clk
		.peripherals_bridge_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // peripherals_bridge_reset_reset_bridge_in_reset.reset
		.peripherals_bridge_m0_address                        (peripherals_bridge_m0_address),                             //                          peripherals_bridge_m0.address
		.peripherals_bridge_m0_waitrequest                    (peripherals_bridge_m0_waitrequest),                         //                                               .waitrequest
		.peripherals_bridge_m0_burstcount                     (peripherals_bridge_m0_burstcount),                          //                                               .burstcount
		.peripherals_bridge_m0_byteenable                     (peripherals_bridge_m0_byteenable),                          //                                               .byteenable
		.peripherals_bridge_m0_read                           (peripherals_bridge_m0_read),                                //                                               .read
		.peripherals_bridge_m0_readdata                       (peripherals_bridge_m0_readdata),                            //                                               .readdata
		.peripherals_bridge_m0_readdatavalid                  (peripherals_bridge_m0_readdatavalid),                       //                                               .readdatavalid
		.peripherals_bridge_m0_write                          (peripherals_bridge_m0_write),                               //                                               .write
		.peripherals_bridge_m0_writedata                      (peripherals_bridge_m0_writedata),                           //                                               .writedata
		.peripherals_bridge_m0_debugaccess                    (peripherals_bridge_m0_debugaccess),                         //                                               .debugaccess
		.epcs_spi_spi_control_port_address                    (mm_interconnect_1_epcs_spi_spi_control_port_address),       //                      epcs_spi_spi_control_port.address
		.epcs_spi_spi_control_port_write                      (mm_interconnect_1_epcs_spi_spi_control_port_write),         //                                               .write
		.epcs_spi_spi_control_port_read                       (mm_interconnect_1_epcs_spi_spi_control_port_read),          //                                               .read
		.epcs_spi_spi_control_port_readdata                   (mm_interconnect_1_epcs_spi_spi_control_port_readdata),      //                                               .readdata
		.epcs_spi_spi_control_port_writedata                  (mm_interconnect_1_epcs_spi_spi_control_port_writedata),     //                                               .writedata
		.epcs_spi_spi_control_port_chipselect                 (mm_interconnect_1_epcs_spi_spi_control_port_chipselect),    //                                               .chipselect
		.gpio_0_s1_address                                    (mm_interconnect_1_gpio_0_s1_address),                       //                                      gpio_0_s1.address
		.gpio_0_s1_write                                      (mm_interconnect_1_gpio_0_s1_write),                         //                                               .write
		.gpio_0_s1_readdata                                   (mm_interconnect_1_gpio_0_s1_readdata),                      //                                               .readdata
		.gpio_0_s1_writedata                                  (mm_interconnect_1_gpio_0_s1_writedata),                     //                                               .writedata
		.gpio_0_s1_chipselect                                 (mm_interconnect_1_gpio_0_s1_chipselect),                    //                                               .chipselect
		.jtag_uart_avalon_jtag_slave_address                  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                    jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                               .write
		.jtag_uart_avalon_jtag_slave_read                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                               .read
		.jtag_uart_avalon_jtag_slave_readdata                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                               .readdata
		.jtag_uart_avalon_jtag_slave_writedata                (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                               .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                               .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect               (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                               .chipselect
		.led_s1_address                                       (mm_interconnect_1_led_s1_address),                          //                                         led_s1.address
		.led_s1_write                                         (mm_interconnect_1_led_s1_write),                            //                                               .write
		.led_s1_readdata                                      (mm_interconnect_1_led_s1_readdata),                         //                                               .readdata
		.led_s1_writedata                                     (mm_interconnect_1_led_s1_writedata),                        //                                               .writedata
		.led_s1_chipselect                                    (mm_interconnect_1_led_s1_chipselect),                       //                                               .chipselect
		.sysid_control_slave_address                          (mm_interconnect_1_sysid_control_slave_address),             //                            sysid_control_slave.address
		.sysid_control_slave_readdata                         (mm_interconnect_1_sysid_control_slave_readdata),            //                                               .readdata
		.systimer_s1_address                                  (mm_interconnect_1_systimer_s1_address),                     //                                    systimer_s1.address
		.systimer_s1_write                                    (mm_interconnect_1_systimer_s1_write),                       //                                               .write
		.systimer_s1_readdata                                 (mm_interconnect_1_systimer_s1_readdata),                    //                                               .readdata
		.systimer_s1_writedata                                (mm_interconnect_1_systimer_s1_writedata),                   //                                               .writedata
		.systimer_s1_chipselect                               (mm_interconnect_1_systimer_s1_chipselect)                   //                                               .chipselect
	);

	cq_viola_irq_mapper irq_mapper (
		.clk           (core_clk),                       //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_e_d_irq_irq)               //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (core_clk),                           //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (peri_clk),                           //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
